* /home/aparna/TBC/Microelectronic_Circuits_:_Theory_And_Applications/CH2/EX2.4/example_2.4/example_2.4.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Wed Aug 26 12:39:35 2015

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
D1  out GND DIODE		
v1  Net-_R1-Pad2_ GND 5V		
R1  out Net-_R1-Pad2_ 1000		

.end
