* EESchema Netlist Version 1.1 (Spice format) creation date: Monday 27 May 2013 03:30:53 PM IST

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

*Sheet Name:/
U1  4 1 VPLOT8_1		
U2  4 3 IPLOT		
R1  1 0 .5k		
v1  4 0 10		
D1  3 1 DIODE		

.end
