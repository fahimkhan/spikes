* eeschema netlist version 1.1 (spice format) creation date: monday 27 may 2013 03:30:53 pm ist

* Plotting option vplot8_1
V_u2 4 3 0
r1  1 0 .5k
v1  4 0 10
d1  3 1 diode

.dc  v1 0e-00 10e-00 100e-03
.plot v(4) v(1) 
.plot i(V_u2)
.end
